module baud_rate_generator (
    input PCLK,             
    input PRESETn,                       
    input spiswai,          
    input [1:0]  spi_mode,         
    input [2:0]  spr,              
    input [2:0]  sppr,                
    input cpol,           
    input  cphase,
    input  ss,            

    output reg sclk,             
    output BaudRateDivisor,  
    output reg   flag_low,         
    output reg   flag_high,        
    output reg   flags_low,        
    output reg   flags_high        
);

reg [11:0] count;
reg pre_sclk = 0;

wire r_mode;
wire w_mode;
wire w1;
wire w2;


assign BaudRateDivisor = ( (sppr + 1 ) * 2^(spr+1) );




assign r_mode = (spi_mode == 2'b00);
assign w_mode = (spi_mode == 2'b01);
assign w1 = ( r_mode || w_mode);
assign w2 = ( w1 && ~ss && ~spiswai);

always@(posedge PCLK  or negedge PRESETn) 
begin
	if(!PRESETn) 
		begin
			count <= 12'b0;
		end
	else if (w2) 
		begin
			if(count == ( BaudRateDivisor -1'b1))
				begin
					count <=12'b0;
				end
			else
				begin
					count <= count +1'b1;
				end
		end
end


always@(posedge PCLK  or negedge PRESETn)
begin
if(!PRESETn) 
		begin
			count <= 12'b0;
		end
	else if (w2) 
		begin
			if(count == ( BaudRateDivisor -1'b1))
				begin
					sclk <= ~sclk;
				end
			else
				begin
					sclk <= sclk;
				end
		end
end

endmodule


